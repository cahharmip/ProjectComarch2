/*
file : Register
By   : Sorapol  Sroysuwan 5610503990
	   Jackthip Phureesatian 5610500966
Date : 9/5/2558
*/

module register (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n,  // Asynchronous reset active low
	
);



endmodule